library ieee;
use ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity ROMModule is
	port(
		IR : in std_logic_vector(15 downto 0);
		clk: in std_logic
	);
end entity ROMModule;

architecture ROMModuleWorkFlow of ROMModule is 
	component PLA 
		PORT(	
			IR    : in std_logic_vector (15 downto 0) ;	
			MPC   : in std_logic_vector(6 downto 0);
   			output: out std_logic_vector (6 downto 0)
		);
	end component;

	component ROM
		port(
			address   : in std_logic_vector(6 downto 0);
			dataOut   : out std_logic_vector(19 downto 0)
		);
	end component;

	component mPCInrementor
		port(
			input : in  std_logic_vector(6 downto 0);
			output: out std_logic_vector(6 downto 0)
		);
	end component;

	signal mPC           : std_logic_vector(6 downto 0);
	signal ROMout        : std_logic_vector(19 downto 0);
	signal PLAOut        : std_logic_vector(6 downto 0);
	signal IncrementedmPC: std_logic_vector(6 downto 0);
	
begin
	ROMX: ROM port map(mPC, ROMout);
	
	PLAX: PLA port map(IR, mPC, PLAOut);
	
	mPCInrementorX: mPCInrementor port map(mPC, IncrementedmPC);
	
	mPC <= PLAOut when (ROMout(10 downto 7) = "1001") and rising_edge(clk) 
	else  mPC or "00000"&IR(8)&"0" when (ROMout(10 downto 7) = "1010") and rising_edge(clk) and mPC(6) = '1' and IR(8) = '1' 
	else  mPC or "00000"&IR(2)&"0" when (ROMout(10 downto 7) = "1010") and rising_edge(clk) and mPC(6) = '0' and IR(2) = '1' 
	else IncrementedmPC when rising_edge(clk) ;

end architecture ROMModuleWorkFlow;