LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY my_adder IS
	PORT (a,b,cin,e: IN  std_logic;
		  s, cout : OUT std_logic );
END my_adder;

ARCHITECTURE a_my_adder OF my_adder IS
	BEGIN
		PROCESS ( a ,b , cin)
			BEGIN 
			IF (e='0')
			Then
				s <= a XOR b XOR cin;
				else
				s<=a;
				end if
				cout <= (a AND b) OR (cin AND (a XOR b));
		END PROCESS;
END a_my_adder;
